`ifndef CLK_IF__SV
`define CLK_IF__SV

interface clk_if();
   logic clk;
endinterface

`endif
