`ifndef A__SV
`define A__SV
class A extends uvm_component;
   `uvm_component_utils(A)

   function new(string name, uvm_component parent);
      super.new(name, parent);
   endfunction

   extern function void build_phase(uvm_phase phase);
   extern virtual  task post_shutdown_phase(uvm_phase phase);
   extern virtual  task run_phase(uvm_phase phase);
endclass

function void A::build_phase(uvm_phase phase);
   super.build_phase(phase);
endfunction

task A::post_shutdown_phase(uvm_phase phase);
   phase.raise_objection(this);
   `uvm_info("A", "post shutdown phase start", UVM_LOW)
   #300;
   `uvm_info("A", "post shutdown phase end", UVM_LOW)
   phase.drop_objection(this);
endtask

task A::run_phase(uvm_phase phase);
   phase.raise_objection(this);
   `uvm_info("A", "run phase start", UVM_LOW)
   #200;
   `uvm_info("A", "run phase end", UVM_LOW)
   phase.drop_objection(this);
endtask

`endif
